module main

import os
import flag
import time

// source https://github.com/enorsu/resource-pack-renamer.git
// feel free to distribute and modify

fn stat(current int, max int) string {
	return '[${current}/${max}] '
}

fn generate_summary(duration i64, total int, proc int) []string {
	return [
		'',
		'SUMMARY:',
		'Processed ${proc} out of the total ${total} files',
		'Process took ${duration}ms',
	]
}

// renaming function
fn rename(blacklist []string, mut files []string, path string) (i64, int, int) {
	// woooo profiling
	sw := time.new_stopwatch()

	// counter variable
	mut i := 0

	// processed files counter
	mut processed_count := 0

	for mut file in files {
		// increment by one
		i = i + 1

		oldfile := file
		// loop through the blacklisted chars
		for item in blacklist {
			// remove char
			file = file.replace(item, '')
		}
		// check if they are equal, so we don't waste no memory
		if oldfile != file {
			// rename(move) the old file
			os.mv('${path}/${oldfile}', '${path}/${file}') or {}

			// print information
			println(stat(i, files.len) + oldfile + ' -> ' + file)
			i += 1
		} else {
			// nothing to do
			println('${stat(i, files.len)}nothing to do')
		}
	}
	return sw.elapsed().milliseconds(), files.len, processed_count
}

fn main() {
	// define blacklisted letters
	mut blacklist := ['[', ']', '(', ')', '!', '§', '¡', '&']

	// initialize flag(argument) parser
	mut fp := flag.new_flag_parser(os.args)

	// set version(s)
	fp.application('resourcepackrenamer')
	fp.version('0.0.1')
	fp.description('rename my packs for me')

	// argument(s)
	path := fp.string('path', `p`, 'none', 'path for processing')

	help := fp.bool('help', `h`, false, 'help')

	if help {
		info := {
			'--help, -h':     'display this'
			'--path, -p':     'set path(required)'
			'--override, -o': 'override list of chars'
		}
		for key, val in info {
			println('${key}     ${val}')
		}
		return
	}
	override := fp.string('override', `o`, 'none', 'override')

	// if user didn't provide a path; return
	if path == 'none' {
		println('a file path is required.')
		println('--help for help')
		return
	}
	// override, overrides the blacklist with a string provided by the user
	if override != 'none' {
		blacklist = override.split('')
	}
	// loop through all the files in the provided location
	mut files := os.ls(path) or { [] }

	duration, total, count := rename(blacklist, mut files, path)
	for item in generate_summary(duration, total, count) {
		println(item)
		println('-'.repeat(item.len))

	}
}
